 `timescale 1ps / 1ps

 module top_module;
   
    reg clk;
    always #5 clk <= ~clk;
    initial 
    begin
        clk = 1'b0;
    end

    dut test(
        .clk(clk));


 endmodule